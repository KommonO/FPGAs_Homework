//Module for the one shot 
module oneshot();



endmodule
