library verilog;
use verilog.vl_types.all;
entity spi_mux_tb is
end spi_mux_tb;
