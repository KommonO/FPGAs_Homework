library verilog;
use verilog.vl_types.all;
entity debounce_tb is
end debounce_tb;
