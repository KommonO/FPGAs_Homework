//Need to create a module for the mux seen in the bottom of the spi wrapper class
//Inputs are 
module spi_mux(input mem_cap, mem_type, man_id, output mux_out);

parameter FFINPUT = 8'hFF;

always @* begin
  


end  //end always @*


endmodule
