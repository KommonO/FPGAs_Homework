//Module to debounce the circuit for the  FPGA board
module debounce();




endmodule 
