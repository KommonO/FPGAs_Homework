//SPI Master for the ST MicroM25P16 Serial Flash
`default_nettype none

module rdid(
  input wire spimiso,
  input wire clk,
  input wire rst,
  input wire get_rdid,
  output reg spisck,
  output wire spimosi,
  output reg prom_cs_n
);

  reg [2:0] current_state, next_state;
  reg [2:0] send_count;
  reg [4:0] get_count;
  reg enable_get_count, enable_send_count;
  reg assert_prom_cs_n;
  wire [7:0] man_id, mem_type, mem_cap;
  reg [23:0] read_data;

  localparam [2:0] SEND_COUNT_MAX = 3'h7;
  localparam [4:0] GET_COUNT_MAX = 5'h18; 
  localparam [7:0] RDID_CMD = 8'h9F; 
  localparam [2:0] IDLE = 3'd0,
    ASSERT_CS=3'd1,
    SEND_INSTRUCTION = 3'd2,
    GET_DATA = 3'd3,
    DEASSERT_CS = 3'd4;
  assign man_id = read_data[23:16];
  assign mem_type = read_data[15:8];
  assign mem_cap = read_data[7:0];

  always @* begin
  //Defaults
  next_state = IDLE;
  enable_send_count = 1'b0;
  enable_get_count = 1'b0;
  assert_prom_cs_n = 1'b0;
  case(current_state)
    //Remain in idle until told to get do RDID
    IDLE: begin
      if (get_rdid)
         next_state = ASSERT_CS;
    end

    ASSERT_CS: begin
      next_state = SEND_INSTRUCTION;
      assert_prom_cs_n = 1'b1;
    end


    //Provide clocks to send the instructions
    SEND_INSTRUCTION: begin
      enable_send_count = 1'b1;
      assert_prom_cs_n = 1'b1; 
      if(send_count == 0)
        next_state = GET_DATA;
      else
        next_state = SEND_INSTRUCTION;
    end

    GET_DATA: begin
      enable_get_count = 1'b1;
      assert_prom_cs_n = 1'b1;
      if(get_count == 0)
        next_state = DEASSERT_CS;
      else
        next_state = GET_DATA;
    end
   

    DEASSERT_CS: begin
      next_state = IDLE;
    end
  endcase
  end
  
  //Need a register so the chip doesnt glitch
  always @(posedge clk or posedge rst) begin
    if(rst)
      prom_cs_n <= 1'b1;
    else if (assert_prom_cs_n)
      prom_cs_n <= 1'b0;
    else
      prom_cs_n <= 1'b1; 
  end
   
  //Current State gets next state at the positive edge of the clock
  always @(posedge clk or posedge rst) begin
    if(rst)
      current_state <= IDLE;
    else
      current_state <= next_state;
  end

  //maintain a count of the spisck's we've provided sending
  always @ (posedge clk or posedge rst) begin
    if(rst)
      send_count <= SEND_COUNT_MAX;
    //rst counter every time we're asked to get the ID again
    else if (get_rdid)
      send_count <= SEND_COUNT_MAX;
    else if (enable_send_count && spisck)
      send_count <= send_count - 1'b1;
  end
  
  //maintain a count of the spisck's we've provided getting
  always @ (posedge clk or posedge rst) begin
    if(rst)
      get_count <= GET_COUNT_MAX;
    else if (get_rdid)
      get_count <= GET_COUNT_MAX;
    else if (enable_get_count && spisck)
      get_count <= get_count - 1'b1; 
  end

  //Collect read_data
  always @(posedge spisck or posedge rst) begin
    if(rst)
      read_data <= 24'b0;
    else 
      read_data[get_count] <= spimiso;
  end

  //Toggle spi_sck need a register so the clock doesnt glitch
  always @ (posedge clk or posedge rst) begin
    if(rst)
      spisck <= 1'b0;
    else if (enable_send_count || enable_get_count)
      spisck <= !spisck;
    else if (get_rdid)
      spisck <= 1'b0;
  end
  
  assign spimosi = RDID_CMD[send_count];
  
  //synopsys_translate off
  reg [250:0] ASCII_current_state, ASCII_next_state; 
  always@* begin
    case(current_state)
      IDLE:ASCII_current_state = "IDLE";
      ASSERT_CS: ASCII_current_state = "ASSERT_CS";
      SEND_INSTRUCTION: ASCII_current_state = "SEND_INSTRUCTION";
      GET_DATA: ASCII_current_state = "GET_DATA";
      DEASSERT_CS: ASCII_current_state = "DEASSERT_CS";
    endcase
  end
  always@* begin
    case(next_state)
      IDLE:ASCII_next_state = "IDLE";
      ASSERT_CS: ASCII_next_state = "ASSERT_CS";
      SEND_INSTRUCTION: ASCII_next_state = "SEND_INSTRUCTION";
      GET_DATA: ASCII_next_state = "GET_DATA";
      DEASSERT_CS: ASCII_next_state = "DEASSERT_CS";
    endcase
  end










endmodule 